`default_nettype none
`include "common_params.h"
`include "common_params_in_fetch_phase.h"

module fetch_phase_displacement (
);
endmodule

`default_nettype wire
